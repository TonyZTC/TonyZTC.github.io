Voltage Divider - Sine
.model Dbreak D Is=1e-16 Rs=0 N=1 TT=0 Cjo=0pF
vin 1 0 sin (0.0V 2.0V 60) ac 1.0 dc 0.0
d1 1 2 Dbreak
r1 2 0 1.0k
.control
tran 0.1ms 30ms
plot v(1) v(2)
.endc
.end
