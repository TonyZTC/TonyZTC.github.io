Voltage Divider - DC
.model Dbreak D Is=1e-16 Rs=0 N=1 TT=0 Cjo=0pF
.DC vin -2 2 0.01
vin 1 0
d1 1 2 Dbreak
r1 2 0 1.0k
.plot DC v(2) 
.end
